`ifndef __JVS_MEMORY_TB_SV__
 `define __JVS_MEMORY_TB_SV__
`include "uvm_macros.svh"
import uvm_pkg::*;
import jvs_pkg::*;

module jvs_memory_tb();
   initial begin
      run_test();
    end
endmodule

`endif
